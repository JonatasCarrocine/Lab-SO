module aluControl(
    input [1:0] aluOp,
    input [5:0] funct,
    output reg [3:0] alu_control
);
    always @(*) begin
        case (aluOp)
            2'b00: alu_control = 4'b0010; // LW/SW/ADDI → ADD
            2'b01: alu_control = 4'b0110; // BEQ → SUB
            2'b10: begin // Tipo R
                case (funct)
                    6'b100000: alu_control = 4'b0010; // ADD
                    6'b100010: alu_control = 4'b0110; // SUB
                    6'b100100: alu_control = 4'b0000; // AND
                    6'b100101: alu_control = 4'b0001; // OR
                    6'b101010: alu_control = 4'b0111; // SLT
                    6'b100111: alu_control = 4'b1100; // NOR
                    default:   alu_control = 4'b0000; // NOP
                endcase
            end
            default: alu_control = 4'b0000;
        endcase
    end
endmodule