module memInstrucao (endInstr, pcInstr, posMem, clock);
	parameter SIZE= 500;
	
	input [31:0] endInstr;
	input clock;
	
	output reg [31:0] pcInstr; //reg atualiza em always
	output reg [31:0] posMem; //reg atualiza em always

	
	reg [31:0] mem [SIZE-1:0];
	reg primeiro_ciclo = 1;
	
	initial
	begin
		//mem[0] = 32'b001100_00000_01000_0000000000000101;// addi 5
		//mem[1] = 32'b001100_00000_01001_0000000000000111;// addi 7
		//mem[2] = 32'b000000_01000_01001_01010_00000_100000;// add
		//mem[3] = 32'b001100_01010_00100_0000000000000000;   //addi $a0, $t2, 0
		//mem[4] = 32'b010110_00000_00100_0000000000000000;   //out $a0
		//mem[5] = 32'b011110_00000_00000_0000000000000000;   //halt
		
		//mem[0] = 32'b001101_00000_11011_0000000000000000;// ldi
		//mem[1] = 32'b001101_00000_11100_0000000000100000;// ldi
		//mem[2] = 32'b001101_00000_11101_0000000000101111;// ldi
		//mem[3] = 32'b010010_00000000000000000000001101;// jmp
		////teste
		//mem[4] = 32'b001110_11011_10001_1111111111111111;// str
		//mem[5] = 32'b001100_11011_00001_0000000000000000;// load
		//mem[6] = 32'b011000_00001_11110_00000_00000000000;// move
		//mem[7] = 32'b000001_11101_11101_1111111111111111;// addi
		//mem[8] = 32'b001100_11101_11111_0000000000000000;// load
		//mem[9] = 32'b010011_11111_00000_0000000000000000;// jr
		//mem[10] = 32'b000001_11101_11101_1111111111111111;// addi
		//mem[11] = 32'b001100_11101_11111_0000000000000000;// load
		//mem[12] = 32'b010011_11111_00000_0000000000000000;// jr
		////main
		//mem[13] = 32'b001100_11011_00010_0000000000000000;// load
		//mem[14] = 32'b001101_00000_00011_0000000000000100;// ldi
		//mem[15] = 32'b011000_00011_00010_00000_00000000000;// move
		//mem[16] = 32'b001110_11011_00010_0000000000000000;// str
		//mem[17] = 32'b001100_11011_00100_0000000000000000;// load
		//mem[18] = 32'b011000_00100_10001_00000_00000000000;// move
		//mem[19] = 32'b000001_11011_11011_0000000000000001;// addi
		//mem[20] = 32'b001101_00000_11111_0000000000011000;// ldi
		//mem[21] = 32'b001110_11101_11111_0000000000000000;// str
		//mem[22] = 32'b000001_11101_11101_0000000000000001;// addi
		//mem[23] = 32'b010010_00000000000000000000000100;// jmp
		//mem[24] = 32'b011000_11110_00101_00000_00000000000;// move
		//mem[25] = 32'b000001_11011_11011_1111111111111111;// addi
		//mem[26] = 32'b011000_00101_10001_00000_00000000000;// move
		//mem[27] = 32'b011000_10001_00110_00000_00000000000;// move
		//mem[28] = 32'b010110_00110_00000_0000000000000000;// out
		//mem[29] = 32'b010100_00000000000000000000000000;// nop
		//mem[30] = 32'b010010_00000000000000000000011111;// jmp
		////end
		//mem[31] = 32'b010111_00000000000000000000000000;// halt
		
		
		mem[0] = 32'b001101_00000_11011_0000000000000000;// ldi
		mem[1] = 32'b001101_00000_11100_0000000000100000;// ldi
		mem[2] = 32'b001101_00000_11101_0000000000101111;// ldi
		mem[3] = 32'b010111_00000000000000000000000000;// halt
	end
	
	
	always @(posedge clock) begin
		if(primeiro_ciclo) begin
			pcInstr <= mem[0]; // no primeiro clock, sai 0
			posMem <= 32'b0;
			primeiro_ciclo <= 0;
		end else begin
			pcInstr <= mem[endInstr]; // depois, busca instrução normalmente
			posMem <= endInstr;
		end
	end
endmodule